localparam [2:0] IDLE_S      = 3'b000;
localparam [2:0] ADD_COLOR_S = 3'b001;
localparam [2:0] DISPLAY_S   = 3'b010;
localparam [2:0] DISPLAY2_S  = 3'b011;
localparam [2:0] INPUT_S     = 3'b100;
localparam [2:0] WIN_S       = 3'b101;
localparam [2:0] LOSE_S      = 3'b110;