module timer(
input CLK,
input RST_N
);

endmodule
