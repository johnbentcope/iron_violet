parameter [2:0] CTRL_IDLE_S      = 3'b000;
parameter [2:0] CTRL_ADD_COLOR_S = 3'b001;
parameter [2:0] CTRL_DISPLAY_S   = 3'b010;
parameter [2:0] CTRL_DISPLAY2_S  = 3'b011;
parameter [2:0] CTRL_INPUT_S     = 3'b100;
parameter [2:0] CTRL_WIN_S       = 3'b101;
parameter [2:0] CTRL_LOSE_S      = 3'b110;

parameter [1:0] TIMR_IDLE_S      = 2'b00;
parameter [1:0] TIMR_COUNT_S     = 2'b00;
